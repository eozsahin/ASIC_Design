module test(
       input wire signed [13:0] inputt,
       output wire signed[13:0] outputt
);


assign outputt = inputt;

endmodule